`timescale 1ns / 1ps

module MatrixVecMul_Core #(
    parameter WIDTH = 24,
    parameter Q = 24'd8380417,
    parameter MU = 26'd33587228 // 2^48 / Q for Barrett
)(
    input  wire          clk,
    input  wire          rst_n,

    // --- ���� Rejsam_a �������� (���� A) ---
    input  wire          i_A_valid,
    input  wire [WIDTH-1:0] i_A_data,
    input  wire [7:0]    i_m_idx,     
    input  wire [3:0]    i_j_idx,     
    input  wire [3:0]    i_l_param,   

    // --- s1 RAM ��ȡ�ӿ� ---
    output wire [7:0]    o_s1_addr,   
    output wire [3:0]    o_s1_poly_idx, 
    input  wire [WIDTH-1:0] i_s1_rdata,  

    // --- �ۼ��� RAM �ӿ� ---
    output wire          o_acc_we,
    output wire [7:0]    o_acc_addr,  // ����ַ (Port A)
    output wire [7:0]    o_acc_waddr, // д��ַ (Port B)
    output wire [WIDTH-1:0] o_acc_wdata,
    input  wire [WIDTH-1:0] i_acc_rdata, // ��ȡ��ǰ�ۼ�ֵ

    // --- ���ս����� ---
    output reg           o_res_valid,
    output reg  [WIDTH-1:0] o_res_data,
    output reg  [7:0]    o_res_m_idx
);

    // ============================================================
    // 1. ��ˮ���ӳٶ���
    // ============================================================
    localparam PIPE_DEPTH = 6; 

    // ============================================================
    // 2. ����ͨ· - �׶� 1: s1 ��ȡ��˷�׼��
    // ============================================================
    assign o_s1_poly_idx = i_j_idx; 
    assign o_s1_addr = i_m_idx; 

    reg [WIDTH-1:0] r_A_data_d1;
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) r_A_data_d1 <= 0;
        else r_A_data_d1 <= i_A_data;
    end

    // ============================================================
    // 3. ����ͨ· - �׶� 2: ģ�� (A * s1 % q)
    // ============================================================
    reg [WIDTH-1:0] mul_op_a, mul_op_b;
    (* use_dsp = "yes" *) reg [2*WIDTH-1:0] prod_reg;
    
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            mul_op_a <= 0;
            mul_op_b <= 0;
            prod_reg <= 0;
        end else begin
            mul_op_a <= r_A_data_d1;
            mul_op_b <= i_s1_rdata; 
            prod_reg <= mul_op_a * mul_op_b;
        end
    end

    wire [WIDTH-1:0] barrett_res;
    // Barrett Լ�� (�ӳ�Լ 3 �ģ������ Stage 5 ��Ч)
    Barrett_reduce #( .WIDTH(WIDTH) ) u_barrett (
        .clk(clk),
        .prod(prod_reg),
        .q(Q),
        .mu(MU),
        .res(barrett_res)
    );

    // ============================================================
    // 4. �����ź��ӳ���
    // ============================================================
    reg [7:0] pipe_m_idx [0:PIPE_DEPTH];
    reg [3:0] pipe_j_idx [0:PIPE_DEPTH];
    reg       pipe_valid [0:PIPE_DEPTH];
    reg [3:0] pipe_l_param [0:PIPE_DEPTH];
    
    integer k;
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            for(k=0; k<=PIPE_DEPTH; k=k+1) begin
                pipe_m_idx[k]   <= 8'd0;
                pipe_j_idx[k]   <= 4'd0;
                pipe_valid[k]   <= 1'b0;
                pipe_l_param[k] <= 4'd0;
            end
        end else begin
            pipe_m_idx[0] <= i_m_idx;
            pipe_j_idx[0] <= i_j_idx;
            pipe_valid[0] <= i_A_valid;
            pipe_l_param[0] <= i_l_param;
            
            for(k=0; k<PIPE_DEPTH; k=k+1) begin
                pipe_m_idx[k+1] <= pipe_m_idx[k];
                pipe_j_idx[k+1] <= pipe_j_idx[k];
                pipe_valid[k+1] <= pipe_valid[k];
                pipe_l_param[k+1] <= pipe_l_param[k];
            end
        end
    end

    // ============================================================
    // 5. ����ͨ· - �׶� 3: ��ȡ & �ۼ� (Stage 5)
    // ============================================================
    
    // [�ؼ��޸� 1] ����ַ��ǰ 1 �� (ʹ�� Stage 4 �ĵ�ַ)
    // �������ݻ��� Stage 5 (PIPE_DEPTH-1) ׼����
    assign o_acc_addr = pipe_m_idx[PIPE_DEPTH-2]; 
    
    // �� Stage 5 ���мӷ�����
    // ��ʱ i_acc_rdata ����Ч�� (��Ӧ pipe_m_idx[PIPE_DEPTH-1])
    // ��ʱ barrett_res Ҳ����Ч�� (���� Barrett ������뵽����)
    
    // ����ǵ�һ�� (j=0)������ RAM ���ݣ���ʼֵΪ 0
    wire [WIDTH-1:0] acc_operand;
    assign acc_operand = (pipe_j_idx[PIPE_DEPTH-1] == 4'd0) ? 24'd0 : i_acc_rdata;

    wire [WIDTH-1:0] add_res;
    mod_add #( .WIDTH(WIDTH) ) u_mod_add (
        .a(barrett_res), // ֱ��ʹ�� Barrett ��������ٶ����ӳ�
        .b(acc_operand),
        .q(Q),
        .res(add_res)
    );

    // [�ؼ��޸� 2] ���ӷ�����Ĵ� 1 ��
    // ����д���������� Stage 6��������Դ�� Stage 5 �ļ�����
    reg [WIDTH-1:0] r_final_res;
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) r_final_res <= 0;
        else r_final_res <= add_res;
    end

    // ============================================================
    // 6. д������� (Stage 6)
    // ============================================================
    
    // дʹ�ܺ͵�ַ������ Stage 6
    assign o_acc_we = pipe_valid[PIPE_DEPTH];
    assign o_acc_waddr = pipe_m_idx[PIPE_DEPTH]; 
    
    // [�ؼ��޸� 3] д����ʹ�üĴ��Ľ��
    assign o_acc_wdata = r_final_res;

    // ��������߼�
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            o_res_valid <= 0;
            o_res_data <= 0;
            o_res_m_idx <= 0;
        end else begin
            if (pipe_valid[PIPE_DEPTH] && (pipe_j_idx[PIPE_DEPTH] == pipe_l_param[PIPE_DEPTH] - 1)) begin
                o_res_valid <= 1'b1;
                o_res_data  <= r_final_res; // ���ҲҪ�üĴ���ֵ
                o_res_m_idx <= pipe_m_idx[PIPE_DEPTH];
            end else begin
                o_res_valid <= 1'b0;
            end
        end
    end

endmodule