`timescale 1ns / 1ps

module Power2Round #(
    parameter WIDTH = 24
)(
    input  wire             clk,
    input  wire             rst_n,
    
    // --- �����ź� ---
    input  wire             i_valid, // ����������Ч��־
    output reg              o_valid, // ���������Ч��־
    
    // --- ���ݽӿ� ---
    input  wire [WIDTH-1:0] i_data,  // ����Ԫ�� t
    output reg  [9:0]       o_t1,    // ��� t1 (�޸�Ϊ 10 bits)
    output reg  [12:0]      o_t0     // ��� t0 (�޸�Ϊ 13 bits)
);
    // --- �������� ---
    // T0_CUTOFF = 2^12 = 4096
    localparam [12:0] T0_CUTOFF = 13'd4096;
    // Case 1 ����: 4096 - (-8192) = 12288
    localparam [13:0] CONST_CASE1 = 14'd12288;
    // Case 2 ����: 4096
    localparam [12:0] CONST_CASE2 = 13'd4096;

    // --- �ڲ��ź� ---
    wire [12:0] t0_raw;
    wire [WIDTH-1:0] t1_raw;

    // 1. ���� t mod 2^13 (ֱ�ӽ�ȡ�� 13 λ)
    assign t0_raw = i_data[12:0];
    // 2. ���� floor(t / 2^13) (ֱ������ 13 λ)
    assign t1_raw = i_data >> 13;

    // --- ���߼� ---
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            o_valid <= 1'b0;
            o_t1    <= 10'd0;
            o_t0    <= 13'd0;
        end else begin
            o_valid <= i_valid;
            if (i_valid) begin
                // MATLAB �߼�ӳ��:
                // if (t0_raw > 2^12)
                //    t0 = 2^12 - (t0_raw - 2^13) = 12288 - t0_raw
                //    t1 = t1_raw + 1
                // else
                //    t0 = 2^12 - t0_raw = 4096 - t0_raw
                //    t1 = t1_raw
                
                if (t0_raw > T0_CUTOFF) begin
                    // Case 1: t0_raw > 4096
                    // t1 ���� 1����Ȼ t1_raw �� 24 λ�������ֵ��Ϊ 1023���� 1 ��Ϊ 1024 (��11λ)
                    // ���� Dilithium ģ���£�t1 ���ֻ�� 1023������ֱ�ӽضϸ�ֵ�� 10 bits ���ɡ�
                    o_t1 <= t1_raw[9:0] + 1'b1;
                    
                    // t0 ���������Ϊ 8191���ʺ� 13 bits
                    o_t0 <= CONST_CASE1 - t0_raw;
                end else begin
                    // Case 2: t0_raw <= 4096
                    o_t1 <= t1_raw[9:0];
                    o_t0 <= CONST_CASE2 - t0_raw;
                end
            end
        end
    end

endmodule