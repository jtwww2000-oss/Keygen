`timescale 1ns / 1ps

module matrix_mul_acc (
    input  wire          clk,
    input  wire          rst_n,
    
    // --- �����ź� ---
    input  wire          i_row_start,
    input  wire          i_is_first_col,
    input  wire          i_is_last_col,
    
    // --- Matrix A ���� (��) ---
    input  wire [22:0]   i_a_data,
    input  wire          i_a_valid,
    
    // --- Vector s1 ���� (���� RAM) ---
    output wire [7:0]    o_s1_addr,
    input  wire [23:0]   i_s1_data,
    
    // --- ������ ---
    output reg           o_res_valid,
    output reg  [23:0]   o_res_data,
    output wire          o_res_last,
    output reg           o_busy
);

    // =========================================================================
    // �������� (�� ntt_core ����һ��)
    // =========================================================================
    localparam [23:0] Q = 24'd8380417;
    localparam [25:0] MU = 26'd33587228; // Barrett Constant for Q

    localparam S_IDLE      = 3'd0;
    localparam S_CALC      = 3'd1;
    localparam S_DUMP_INIT = 3'd2;
    localparam S_DUMP      = 3'd3;
    localparam S_DONE      = 3'd4;
    
    reg [2:0] state;

    // =========================================================================
    // �ڲ��ź�
    // =========================================================================
    reg [8:0] cnt;
    
    // FIFO
    wire        fifo_empty;
    wire        fifo_rd_en;
    wire [22:0] fifo_a_out;
    
    // �˷��� (DSP + Barrett)
    (* use_dsp = "yes" *) reg [47:0] prod_reg; // 23bit * 24bit -> 47bit
    wire [23:0] mul_res;
    
    // �ӷ���
    wire [23:0] add_res;
    
    // �ۼ��� RAM
    reg  [7:0]  acc_addr_rd;
    reg  [7:0]  acc_addr_wr;
    reg         acc_we;
    reg  [23:0] acc_wdata;
    wire [23:0] acc_rdata;
    
    // ��ˮ�߿���
    reg         pipe_valid_s1; 
    reg         pipe_valid_mult;
    reg         pipe_is_first_col; 
    reg [7:0]   pipe_addr_stage1;
    reg [7:0]   pipe_addr_stage2;

    // =========================================================================
    // 1. ���� FIFO
    // =========================================================================
    simple_fifo #( .WIDTH(23), .DEPTH(16) ) u_a_fifo (
        .clk(clk), .rst_n(rst_n),
        .we(i_a_valid), .din(i_a_data),
        .re(fifo_rd_en), .dout(fifo_a_out),
        .empty(fifo_empty), .full()
    );

    // =========================================================================
    // 2. �������߼�
    // =========================================================================
    assign fifo_rd_en = (state == S_CALC) && (!fifo_empty);
    assign o_s1_addr = cnt[7:0];

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= S_IDLE;
            cnt <= 0;
            o_busy <= 0;
            pipe_valid_s1 <= 0;
            pipe_valid_mult <= 0;
            pipe_is_first_col <= 0;
            acc_we <= 0;
        end else begin
            acc_we <= 0;
            
            case (state)
                S_IDLE: begin
                    o_busy <= 0;
                    if (i_row_start) begin
                        state <= S_CALC;
                        cnt <= 0;
                        o_busy <= 1;
                    end
                end

                S_CALC: begin
                    // --- Stage 0: Request ---
                    if (!fifo_empty) begin
                        pipe_valid_s1 <= 1;
                        pipe_is_first_col <= i_is_first_col;
                        pipe_addr_stage1 <= cnt[7:0];
                        
                        if (cnt == 255) cnt <= 0;
                        else cnt <= cnt + 1;
                    end else begin
                        pipe_valid_s1 <= 0;
                    end

                    // --- Stage 1: Multiply Input Latch ---
                    if (pipe_valid_s1) begin
                        // ׼���˷�����: A * s1
                        prod_reg <= fifo_a_out * i_s1_data; 
                        
                        pipe_valid_mult <= 1;
                        pipe_addr_stage2 <= pipe_addr_stage1;
                        acc_addr_rd <= pipe_addr_stage1; 
                    end else begin
                        pipe_valid_mult <= 0;
                    end

                    // --- Stage 2: Add & Write Back ---
                    // Barrett Լ����Ľ���� mul_res �� (����߼�/�ڲ���ˮ)
                    if (pipe_valid_mult) begin
                        acc_we <= 1;
                        acc_addr_wr <= pipe_addr_stage2;
                        
                        if (pipe_is_first_col) begin
                            acc_wdata <= mul_res; // ��һ��ֱ�Ӹ���
                        end else begin
                            acc_wdata <= add_res; // �������ۼ�
                        end
                        
                        // ����Ƿ���һ�е����һ������
                        if (pipe_addr_stage2 == 255 && i_is_last_col) begin
                            state <= S_DUMP_INIT;
                        end
                    end
                end

                S_DUMP_INIT: begin
                    cnt <= 0;
                    acc_we <= 0;
                    acc_addr_rd <= 0;
                    state <= S_DUMP;
                end

                S_DUMP: begin
                    if (cnt < 256) begin
                        o_res_valid <= (cnt > 0); 
                        o_res_data  <= acc_rdata;
                        if (cnt < 255) acc_addr_rd <= cnt[7:0] + 1;
                        cnt <= cnt + 1;
                    end else begin
                        o_res_valid <= 1;
                        o_res_data  <= acc_rdata;
                        state <= S_DONE;
                    end
                end
                
                S_DONE: begin
                    o_res_valid <= 0;
                    o_busy <= 0;
                    state <= S_IDLE;
                end
            endcase
        end
    end
    
    assign o_res_last = (state == S_DONE);

    // =========================================================================
    // 3. ���㵥Ԫʵ���� (FIXED)
    // =========================================================================
    
    // [FIX] ʹ�� Barrett_reduce ��� Montgomery_mul���� ntt_core һ��
    Barrett_reduce #( .WIDTH(24) ) u_barrett (
        .clk(clk),
        .prod(prod_reg),
        .q(Q),
        .mu(MU),
        .res(mul_res) // �˷���� A*s1 mod Q
    );
    
    // [FIX] ���� mod_add �ӿ�
    mod_add #( .WIDTH(24) ) u_add (
        .a(acc_rdata),
        .b(mul_res),
        .q(Q),         // ����ȱ�� Q ����
        .res(add_res)  // �����˿��� c -> res
    );

    // =========================================================================
    // 4. �ۼ��� RAM
    // =========================================================================
    tdpram_24x256_internal u_acc_ram (
        .clk(clk),
        .we_a(1'b0), .addr_a(acc_addr_rd), .din_a(24'd0), .dout_a(acc_rdata),
        .we_b(acc_we), .addr_b(acc_addr_wr), .din_b(acc_wdata), .dout_b()
    );

endmodule

// Helper modules (FIFO & RAM) kept same as before...
module simple_fifo #(parameter WIDTH=23, DEPTH=16) (
    input wire clk, rst_n, we, input wire [WIDTH-1:0] din,
    input wire re, output wire [WIDTH-1:0] dout, output wire empty, output wire full
);
    reg [WIDTH-1:0] mem [0:DEPTH-1];
    reg [4:0] wptr, rptr;
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin wptr<=0; rptr<=0; end
        else begin
            if (we && !full) begin mem[wptr[3:0]]<=din; wptr<=wptr+1; end
            if (re && !empty) rptr<=rptr+1;
        end
    end
    assign dout = mem[rptr[3:0]];
    assign empty = (wptr == rptr);
    assign full  = (wptr[3:0] == rptr[3:0]) && (wptr[4] != rptr[4]);
endmodule

module tdpram_24x256_internal (
    input wire clk,
    input wire we_a, input wire [7:0] addr_a, input wire [23:0] din_a, output reg [23:0] dout_a,
    input wire we_b, input wire [7:0] addr_b, input wire [23:0] din_b, output reg [23:0] dout_b
);
    reg [23:0] ram [0:255];
    integer i;
    initial begin for(i=0; i<256; i=i+1) ram[i] = 0; end
    always @(posedge clk) begin if (we_a) ram[addr_a] <= din_a; dout_a <= ram[addr_a]; end
    always @(posedge clk) begin if (we_b) ram[addr_b] <= din_b; dout_b <= ram[addr_b]; end
endmodule