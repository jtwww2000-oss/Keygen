`timescale 1ns / 1ps

module pk_packer (
    input  wire          clk,
    input  wire          rst_n,
    
    // --- ���� ---
    input  wire          start_pack, // �� rho ׼����ʱ����
    
    // --- �������� ---
    input  wire [255:0]  rho,
    input  wire          t1_valid,
    input  wire [9:0]    t1_data,
    
    // --- �����λ��Կ ---
    // Max size for Dilithium5: 256 (rho) + 8*256*10 (t1) = 20736 bits
    output reg [20735:0] o_pk_bus,  
    output reg           o_pk_done    // ���������ݴ�����ʱ����
);

    // ָ�룬ָʾ��ǰд���λ��
    // ���λ�� 20736����Ҫ 15 bits (2^15 = 32768)
    reg [14:0] write_ptr;
    
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            o_pk_bus   <= 0;
            write_ptr  <= 0;
            o_pk_done  <= 0;
        end else begin
            // ����ʱ���� rho ���� 256 λ
            if (start_pack) begin
                o_pk_bus[255:0] <= rho;
                write_ptr       <= 256;
                o_pk_done       <= 0;
                // �����λ������ (��ѡ)
                o_pk_bus[20735:256] <= 0;
            end
            
            // �� t1 ��Чʱ��ƴ�ӵ���ǰָ��λ��
            if (t1_valid) begin
                // Verilog �Ķ�̬λ��Ƭ�﷨: [base +: width]
                // �� 10-bit t1 д�뵱ǰ write_ptr ��ʼ�� 10 λ
                o_pk_bus[write_ptr +: 10] <= t1_data;
                
                // ָ�벽��
                write_ptr <= write_ptr + 10;
            end
            
            // �жϽ������� (��������ⲿ��λ����һ�� start �������
            // ��������Ը��� write_ptr ��ֵ���ж� done)
            // Dilithium2: 256 + 4*256*10 = 10496
            // Dilithium3: 256 + 6*256*10 = 15616
            // Dilithium5: 256 + 8*256*10 = 20736
            // ����������һ���򵥵��߼�������ںܳ�һ��ʱ��û�� valid �źţ����� KeyGen ����ˣ�
            // �ϲ�ģ���������̡���ģ�������"�ۼ�"��
            // Ϊ�˷�����ԣ����ǿ��Լ���ض��� write_ptr ֵ���� done��
            // ��Ϊ��ͨ���ԣ������� KeyGen �� done �ź�ֱ�������ⲿ�۲졣
        end
    end

endmodule